*  Generated for: PrimeSim
*  Design library name: Dynamic_CP
*  Design cell name: Dynamic_CP_Circuit_tb
*  Design view name: schematic
.lib 'saed32nm.lib' TT

*Custom Compiler Version S-2021.09
*Wed Feb 23 21:50:30 2022

.global gnd!
********************************************************************************
* Library          : Dynamic_CP
* Cell             : Dynamic_CP_Circuit
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt dynamic_cp_circuit clk1 clk2 gnd_1 out vdd
xm16 clk2 vdd net70 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm11 clk1 vdd net50 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm6 clk2 vdd net30 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm0 clk1 vdd net101 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm23 net84 out net92 net92 p105 w=0.1u l=0.03u nf=1 m=1
xm22 net92 net84 out net92 p105 w=0.1u l=0.03u nf=1 m=1
xm21 net84 out out net92 p105 w=0.1u l=0.03u nf=1 m=1
xm20 net72 net84 net80 net80 p105 w=0.1u l=0.03u nf=1 m=1
xm19 net80 net72 net84 net80 p105 w=0.1u l=0.03u nf=1 m=1
xm18 net72 net70 net84 net80 p105 w=0.1u l=0.03u nf=1 m=1
xm17 net70 net72 net84 net80 p105 w=0.1u l=0.03u nf=1 m=1
xm15 net52 net72 net60 net60 p105 w=0.1u l=0.03u nf=1 m=1
xm14 net60 net52 net72 net60 p105 w=0.1u l=0.03u nf=1 m=1
xm13 net52 net50 net72 net60 p105 w=0.1u l=0.03u nf=1 m=1
xm12 net50 net52 net72 net60 p105 w=0.1u l=0.03u nf=1 m=1
xm10 net103 net52 net40 net40 p105 w=0.1u l=0.03u nf=1 m=1
xm9 net40 net103 net52 net40 p105 w=0.1u l=0.03u nf=1 m=1
xm8 net103 net30 net52 net40 p105 w=0.1u l=0.03u nf=1 m=1
xm7 net30 net103 net52 net40 p105 w=0.1u l=0.03u nf=1 m=1
xm5 net102 vdd net103 net102 p105 w=0.1u l=0.03u nf=1 m=1
xm4 vdd net103 net102 net102 p105 w=0.1u l=0.03u nf=1 m=1
xm3 vdd net101 net103 net102 p105 w=0.1u l=0.03u nf=1 m=1
xm1 net101 vdd net103 net102 p105 w=0.1u l=0.03u nf=1 m=1
c35 net84 clk2 c=20p
c34 net72 clk1 c=20p
c33 net52 clk2 c=20p
c32 net103 clk1 c=20p
.ends dynamic_cp_circuit

********************************************************************************
* Library          : Dynamic_CP
* Cell             : Dynamic_CP_Circuit_tb
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
xi0 clk1 clk2 gnd! out in dynamic_cp_circuit
v19 clk2 gnd! dc=0 pulse ( 0 'x' 0 0.01u 0.01u 0.25u 0.5u )
v18 clk1 gnd! dc=0 pulse ( 'x' 0 0 0.01u 0.01u 0.25u 0.5u )
c24 out gnd! c=40p
v26 in gnd! dc='x'
r17 out gnd! r=1meg








.tran '1u' '40u' name=tran

.option primesim_remove_probe_prefix = 0
.probe v(*) i(*) level=1
.probe tran v(out)

.temp 25



.option primesim_output=wdf


.option parhier = LOCAL






.end
